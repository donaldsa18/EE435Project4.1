
package states;
typedef enum {GR,YR,RG,RY} state_t;
typedef enum {G,Y,R} light_t;
endpackage